//func
`define addu  6'b100001
`define subu  6'b100011
`define jr    6'b001000
`define slt   6'b101010

//opcode
`define lw   6'b100011
`define lb   6'b100000
`define addi 6'b001000
`define addiu 6'b001001
`define beq  6'b000100
`define sw   6'b101011
`define lui  6'b001111
`define j    6'b000010
`define jal  6'b000011
`define ori  6'b001101